module main
import setuper { setup }

setup(
	name='setuper',
	version='1.0.0',
	repo='https://github.com/v-libs/setuper',
	license='MIT',
	author='snxx',
	email='snxx.lppxx@gmail.com',
	description='Easily create modules'
)
