module setuper

import os

pub fn windows_only() {
	if os.name == 'nt' {
		return args, kwargs
	}

	return func
}
