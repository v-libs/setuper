module setuper

pub fn get_unpatched() {

}

pub fn get_unpatched_class() {

}

pub fn patch_all() {

}

pub fn patch_func() {

}

pub fn get_unpatched_func() {

}