module setuper

import sys
import os
