module setuper
